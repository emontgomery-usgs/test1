netcdf 7751wh {
dimensions:
	time = UNLIMITED ; // (5179 currently)
	depth = xxdepthxx ;
	lon = 1 ;
	lat = 1 ;
variables:
	int time(time) ;
		time:FORTRAN_format = "F10.2" ;
		time:units = "True Julian Day" ;
		time:type = "UNEVEN" ;
		time:epic_code = 624 ;
		time:_FillValue = 0 ;
	int time2(time) ;
		time2:FORTRAN_format = "F10.2" ;
		time2:units = "msec since 0:00 GMT" ;
		time2:type = "UNEVEN" ;
		time2:epic_code = 624 ;
		time2:_FillValue = 0 ;
	float depth(depth) ;
		depth:FORTRAN_format = "F10.2" ;
		depth:units = "m" ;
		depth:type = "EVEN" ;
		depth:epic_code = 3 ;
		depth:long_name = "DEPTH (m)" ;
		depth:blanking_distance = 1.75999999046326 ;
		depth:bin_size = 2. ;
		depth:xducer_offset_from_bottom = 3.33999991416931 ;
		depth:_FillValue = 1.e+35f ;
		depth:NOTE = "Depth values were calculated using Surface.exe output" ;
	float lon(lon) ;
		lon:FORTRAN_format = "f10.4" ;
		lon:units = "degree_east" ;
		lon:type = "EVEN" ;
		lon:epic_code = 502 ;
		lon:name = "LON" ;
		lon:long_name = "LONGITUDE" ;
		lon:generic_name = "lon" ;
		lon:_FillValue = 1.e+35f ;
	float lat(lat) ;
		lat:FORTRAN_format = "F10.2" ;
		lat:units = "degree_north" ;
		lat:type = "EVEN" ;
		lat:epic_code = 500 ;
		lat:name = "LAT" ;
		lat:long_name = "LATITUDE" ;
		lat:generic_name = "lat" ;
		lat:_FillValue = 1.e+35f ;
	float u_1205(time, depth, lat, lon) ;
		u_1205:name = "u" ;
		u_1205:long_name = "Eastward Velocity" ;
		u_1205:generic_name = "u" ;
		u_1205:FORTRAN_format = " " ;
		u_1205:units = "cm/s" ;
		u_1205:epic_code = 1205 ;
		u_1205:sensor_type = "RD Instruments ADCP" ;
		u_1205:sensor_depth = 29.3871691226959 ;
		u_1205:serial_number = 185 ;
		u_1205:minimum = -103.6494f ;
		u_1205:maximum = 109.0786f ;
		u_1205:valid_range = 1000.f, 1000.f ;
		u_1205:_FillValue = 1.e+35f ;
	float v_1206(time, depth, lat, lon) ;
		v_1206:name = "v" ;
		v_1206:long_name = "Northward Velocity" ;
		v_1206:generic_name = "v" ;
		v_1206:FORTRAN_format = " " ;
		v_1206:units = "cm/s" ;
		v_1206:epic_code = 1206 ;
		v_1206:sensor_type = "RD Instruments ADCP" ;
		v_1206:sensor_depth = 29.3871691226959 ;
		v_1206:serial_number = 185 ;
		v_1206:minimum = -104.6426f ;
		v_1206:maximum = 105.0741f ;
		v_1206:valid_range = 1000.f, 1000.f ;
		v_1206:_FillValue = 1.e+35f ;
	float AGC_1202(time, depth, lat, lon) ;
		AGC_1202:name = "AGC" ;
		AGC_1202:long_name = "Average Echo Intensity (AGC)" ;
		AGC_1202:generic_name = "AGC" ;
		AGC_1202:FORTRAN_format = "F5.1" ;
		AGC_1202:units = "counts" ;
		AGC_1202:epic_code = 1202 ;
		AGC_1202:sensor_type = "RD Instruments ADCP" ;
		AGC_1202:sensor_depth = 29.3871691226959 ;
		AGC_1202:serial_number = 185 ;
		AGC_1202:norm_factor = 0.449999988079071 ;
		AGC_1202:NOTE = "normalization to db" ;
		AGC_1202:minimum = 63.75f ;
		AGC_1202:maximum = 215.75f ;
		AGC_1202:valid_range = 50., 255. ;
		AGC_1202:_FillValue = 1.e+35f ;
	float corrl(time, depth, lat, lon) ;
		corrl:name = "PGd" ;
		corrl:long_name = "Percent Good Pings" ;
		corrl:generic_name = "PGd" ;
		corrl:FORTRAN_format = " " ;
		corrl:units = "counts" ;
		corrl:epic_code = 1203 ;
		corrl:sensor_type = "RD Instruments ADCP" ;
		corrl:sensor_depth = 29.3871691226959 ;
		corrl:serial_number = 185 ;
		corrl:minimum = 10.5f ;
		corrl:maximum = 100.f ;
		corrl:valid_range = 0., 100. ;
		corrl:_FillValue = 1.e+35f ;
	float sstrn(time, lat, lon) ;
		sstrn:name = "hght" ;
		sstrn:long_name = "height of sea surface" ;
		sstrn:generic_name = "height" ;
		sstrn:FORTRAN_format = "f10.2" ;
		sstrn:units = "m" ;
		sstrn:epic_code = 18 ;
		sstrn:sensor_depth = 29.3871691226959 ;
		sstrn:minimum = 26.33f ;
		sstrn:maximum = 31.53f ;
		sstrn:serial_number = 185 ;
		sstrn:valid_range = 0.f, 1000.f ;
		sstrn:_FillValue = 1.e+35f ;
		sstrn:NOTE = "height of sea surface relative to transducer head from surface.exe" ;

// global attributes:
		:CREATION_DATE = "15-Feb-2005 15:10:54" ;
		:MOORING = "LA00A5" ;
		:Deployment_date = "09-sep-2004" ;
		:Recovery_date = "09-feb-2005" ;
		:INST_TYPE = "Sontek ADP" ;
		:history = "ASCII files sent to USGS April, 2007. Converted to netcdf using n_rdlacsd.m and n_wrtnc.m" ;
		:firmware_version = 6.7f ;
		:frequency = 500 ;
		:beam_pattern = "convex" ;
		:orientation = "UP" ;
		:beam_angle = 30 ;
		:janus = "4 Beam" ;
		:pings_per_ensemble = 300 ;
		:ADP_serial_number = 251 ;
		:transform = "EARTH" ;
		:DATA_TYPE = "ADCP" ;
		:DATA_SUBTYPE = "MOORED" ;
		:DATA_ORIGIN = "Los Angeles County Sanitation Districts" ;
		:COORD_SYSTEM = "GEOGRAPHIC" ;
		:WATER_MASS = "?" ;
		:POS_CONST = 0 ;
		:DEPTH_CONST = 0 ;
		:WATER_DEPTH = 32.7271690368652 ;
		:DRIFTER = 0 ;
		:VAR_FILL = 1.00000004091848e+35 ;
		:EXPERIMENT = "LACSD Palos Verdes" ;
		:PROJECT = "LACSD" ;
		:DESCRIPT = "A5 ADP" ;
		:longitude = -70.7808 ;
		:latitude = 42.3786 ;
		:DATA_CMNT = "metadata may be wrong" ;
		:FILL_FLAG = 1 ;
		:COMPOSITE = 0 ;
		:VAR_DESC = "u:v:AGC:corr:sstrn" ;
		:DELTA_T = "900" ;
		:start_time = "22-Sep-2004 15:12:30" ;
		:stop_time = "15-Nov-2004 13:42:30" ;
		:magnetic_variation = 13.6 ;
}
