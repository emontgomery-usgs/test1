netcdf 7751wh {
dimensions:
	time = UNLIMITED ; // (5179 currently)
	depth = xxdepthxx ;
	lon = 1 ;
	lat = 1 ;
variables:
	int time(time) ;
		time:FORTRAN_format = "F10.2" ;
		time:units = "True Julian Day" ;
		time:type = "UNEVEN" ;
		time:epic_code = 624 ;
	int time2(time) ;
		time2:FORTRAN_format = "F10.2" ;
		time2:units = "msec since 0:00 GMT" ;
		time2:type = "UNEVEN" ;
		time2:epic_code = 624 ;
	float depth(depth) ;
		depth:FORTRAN_format = "F10.2" ;
		depth:units = "m" ;
		depth:type = "EVEN" ;
		depth:epic_code = 3 ;
		depth:long_name = "DEPTH (m)" ;
		depth:blanking_distance = 1.0 ;
		depth:bin_size = 3. ;
		depth:NOTE = "Depth from LACSD file, line 1" ;
	float lon(lon) ;
		lon:FORTRAN_format = "f10.4" ;
		lon:units = "degree_east" ;
		lon:type = "EVEN" ;
		lon:epic_code = 502 ;
		lon:name = "LON" ;
		lon:long_name = "LONGITUDE" ;
		lon:generic_name = "lon" ;
	float lat(lat) ;
		lat:FORTRAN_format = "F10.2" ;
		lat:units = "degree_north" ;
		lat:type = "EVEN" ;
		lat:epic_code = 500 ;
		lat:name = "LAT" ;
		lat:long_name = "LATITUDE" ;
		lat:generic_name = "lat" ;
	float u_1205(time, depth, lat, lon) ;
		u_1205:name = "u" ;
		u_1205:long_name = "Eastward Velocity" ;
		u_1205:generic_name = "u" ;
		u_1205:FORTRAN_format = " " ;
		u_1205:units = "cm/s" ;
		u_1205:epic_code = 1205 ;
		u_1205:sensor_type = "Sontek ADP" ;
		u_1205:sensor_depth = 65 ;
		u_1205:serial_number = 251 ;
		u_1205:minimum = -103.6494f ;
		u_1205:maximum = 109.0786f ;
		u_1205:valid_range = 1000.f, 1000.f ;
		u_1205:_FillValue = 1.e+35f ;
	float v_1206(time, depth, lat, lon) ;
		v_1206:name = "v" ;
		v_1206:long_name = "Northward Velocity" ;
		v_1206:generic_name = "v" ;
		v_1206:FORTRAN_format = " " ;
		v_1206:units = "cm/s" ;
		v_1206:epic_code = 1206 ;
		v_1206:sensor_type = "Sontek ADP" ;
		v_1206:sensor_depth = 65 ;
		v_1206:serial_number = 251 ;
		v_1206:minimum = -104.6426f ;
		v_1206:maximum = 105.0741f ;
		v_1206:valid_range = 1000.f, 1000.f ;
		v_1206:_FillValue = 1.e+35f ;
	float ampl(time, depth, lat, lon) ;
		ampl:name = "ampl" ;
		ampl:long_name = "4-head averaged Returned transmit signal amplitude (strength)" ;
		ampl:generic_name = "AGC" ;
		ampl:FORTRAN_format = "F5.1" ;
		ampl:units = "counts" ;
		ampl:sensor_type = "Sontek ADP" ;
		ampl:sensor_depth = 65 ;
		ampl:serial_number = 251 ;
		ampl:norm_factor = 1 ;
		ampl:NOTE = "cannot be converted to db; these are in counts" ;
		ampl:minimum = 63.75f ;
		ampl:maximum = 215.75f ;
		ampl:valid_range = 0.f, 255.f ;
		ampl:_FillValue = 1.e+35f ;
	float snr(time, depth, lat, lon) ;
		snr:name = "SNR" ;
		snr:long_name = "4-head averaged Signal-to-noise ratio of the received signal" ;
		snr:generic_name = "SNR" ;
		snr:FORTRAN_format = " " ;
		snr:units = "dB" ;
		snr:sensor_type = "Sontek ADP" ;
		snr:sensor_depth = 65 ;
		snr:serial_number = 251 ;
		snr:minimum = 10.5f ;
		snr:maximum = 100.f ;
		snr:valid_range = 0.f, 100.f ;
		snr:_FillValue = 1.e+35f ;
	float stdcor(time, depth, lat, lon) ;
		stdcor:name = "stdcor" ;
		stdcor:long_name = "4-head averaged Standard Deviation / Correlation of the velocity" ;
		stdcor:sensor_type = "Sontek ADP" ;
		stdcor:generic_name = " stdcor" ;
		stdcor:FORTRAN_format = "f10.2" ;
		stdcor:units = "cm/s" ;
		stdcor:sensor_depth = 65 ;
		stdcor:minimum = 26.33f ;
		stdcor:maximum = 31.53f ;
		stdcor:serial_number = 251 ;
		stdcor:valid_range = 0.f, 50.f ;
		stdcor:_FillValue = 1.e+35f ;

// global attributes:
		:CREATION_DATE = "15-Feb-2005 15:10:54" ;
		:MOORING = "LA00A5" ;
		:Deployment_date = "09-sep-2004" ;
		:Recovery_date = "09-feb-2005" ;
		:INST_TYPE = "Sontek ADP" ;
		:history = "ASCII files sent to USGS April, 2007. Converted to netcdf using n_rdlacsd.m and n_wrtnc.m" ;
		:firmware_version = 6.7f ;
		:frequency = 500 ;
		:beam_pattern = "convex" ;
		:orientation = "UP" ;
		:beam_angle = 30 ;
		:janus = "4 Beam" ;
		:ADP_serial_number = 251 ;
		:transform = "EARTH" ;
		:DATA_TYPE = "ADCP" ;
		:DATA_SUBTYPE = "MOORED" ;
		:DATA_ORIGIN = "Los Angeles County Sanitation Districts" ;
		:COORD_SYSTEM = "GEOGRAPHIC" ;
		:WATER_MASS = "?" ;
		:POS_CONST = 0 ;
		:DEPTH_CONST = 0 ;
		:WATER_DEPTH = 32.7271690368652 ;
		:DRIFTER = 0 ;
		:VAR_FILL = 1.00000004091848e+35 ;
		:EXPERIMENT = "LACSD Palos Verdes" ;
		:PROJECT = "LACSD" ;
		:DESCRIPT = "A5 ADP" ;
		:longitude = -70.7808 ;
		:latitude = 42.3786 ;
		:DATA_CMNT = "metadata from ascii headers- may be incomplete" ;
		:FILL_FLAG = 1 ;
		:COMPOSITE = 0 ;
		:VAR_DESC = "u:v:ampl:snr:stdcor" ;
		:DELTA_T = "900" ;
		:start_time = "22-Sep-2004 15:12:30" ;
		:stop_time = "15-Nov-2004 13:42:30" ;
		:magnetic_variation = 13.6 ;
}
